library verilog;
use verilog.vl_types.all;
entity forwarding is
end forwarding;
