library verilog;
use verilog.vl_types.all;
entity controller is
    port(
        op              : in     vl_logic_vector(5 downto 0);
        funct           : in     vl_logic_vector(5 downto 0);
        zero            : in     vl_logic;
        signext         : out    vl_logic;
        shiftl16        : out    vl_logic;
        memtoreg        : out    vl_logic_vector(1 downto 0);
        memwrite        : out    vl_logic;
        pcsrc           : out    vl_logic;
        alusrc          : out    vl_logic;
        regdst          : out    vl_logic_vector(1 downto 0);
        regwrite        : out    vl_logic;
        jump            : out    vl_logic_vector(1 downto 0);
        alucontrol      : out    vl_logic_vector(2 downto 0);
        jrjump          : out    vl_logic_vector(1 downto 0)
    );
end controller;
